`include "arith.v"

module top (

);
endmodule
